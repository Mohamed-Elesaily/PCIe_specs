module timer (input clk,input [5:0]setTimer,input enableTimer,input resetTimer,output timeOut);

assign timeOut = 1'b0;
endmodule
